// To work with our autograder you MUST be able to get your cpu.v to work
// without making ANY changes to this file.  Refer to Section 4 in the Lab
// 6 handout for more details.




module cpu_autograder_example_tb;
  

reg clk, reset, s, load;
  
reg [15:0] in;
  
wire [15:0] out;
  
wire N,V,Z,w;

  
reg err;

  


cpu DUT(clk,reset,s,load,in,out,N,V,Z,w);

  

initial begin
    
clk = 0; #5;
    
forever begin
      
clk = 1; #5;
      
clk = 0; #5;
    
end
  
end

  
initial begin
    
err = 0;
    
reset = 1; 
s = 0; 
load = 0; 
in = 16'b0;
    
#10;
    
reset = 0; 
    
#10;

    
in = 16'b1101000000000111;
    
load = 1;
    
#10;
    
load = 0;
    
s = 1;
    
#10
    

s = 0;
    @(posedge w); 
// wait for w to go high again
    
#10;
    
if (cpu_autograder_example_tb.DUT.DP.REGFILE.R0 !== 16'h7) begin
      
err = 1;
      
$display("FAILED: MOV R0, #7");
      
$stop;
    
end

    in = 16'b1101000100000010;
    
load = 1;
   
 #10;
    
load = 0;
    
s = 1;
    
#10
    
s = 0;
    
@(posedge w); 
// wait for w to go high again
   
 #10;
    
if (cpu_autograder_example_tb.DUT.DP.REGFILE.R1 !== 16'h2) 
begin
      
err = 1;
      
$display("FAILED: MOV R1, #2");
      
$stop;
    
end

    
in = 16'b1010000101001000;
    
load = 1;
    
#10;
    
load = 0;
    
s = 1;
    
#10
    
s = 0;
   
@(posedge w); // wait for w to go high again
    
#10;
    
if (cpu_autograder_example_tb.DUT.DP.REGFILE.R2 !== 16'h10) 
begin
      
err = 1;
     
 $display("FAILED: ADD R2, R1, R0, LSL#1");
      
$stop;
    
end
    
if (~err) $display("INTERFACE OK");
    
$stop;
  
end
endmodule
